module _XOR(A,B,Y); //XOR gate by using inverter,and,or
input A,B; // declear to input value
output Y;  // declear to see result

assign Y = A ^ B; //assign : ^ is ⊕

endmodule
